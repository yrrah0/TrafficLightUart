library verilog;
use verilog.vl_types.all;
entity txTest_vlg_vec_tst is
end txTest_vlg_vec_tst;
