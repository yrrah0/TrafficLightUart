library verilog;
use verilog.vl_types.all;
entity BaudTest_vlg_vec_tst is
end BaudTest_vlg_vec_tst;
